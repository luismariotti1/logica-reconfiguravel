LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;

ENTITY ConversorCodBinarioGrayGenerateCondicional IS
    PORT (
        entradas : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
        saidas : OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
    );
END ConversorCodBinarioGrayGenerateCondicional;

ARCHITECTURE logic OF ConversorCodBinarioGrayGenerateCondicional IS
BEGIN
    gen : FOR i IN 3 DOWNTO 0 GENERATE
        gen1 : IF i = 3 GENERATE
            saidas(i) <= entradas(i);
        END GENERATE gen1;
        gen2 : IF i /= 3 GENERATE
            saidas(i) <= entradas(i + 1) XOR entradas(i);
        END GENERATE gen2;
    END GENERATE gen;
END logic;