LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;

ENTITY Mux4Por1When8Bits IS
    PORT (
        SELETOR : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
        SAIDA : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
    );

END Mux4Por1When8Bits;

ARCHITECTURE logica OF Mux4Por1When8Bits IS
BEGIN
    SAIDA <= "11000000" WHEN SELETOR = "00" ELSE
        "00110000" WHEN SELETOR = "01" ELSE
        "00001100" WHEN SELETOR = "10" ELSE
        "00000011" WHEN SELETOR = "11";
END logica;